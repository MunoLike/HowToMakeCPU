library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.std_logic_unsigned.all;

